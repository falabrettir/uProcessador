library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity uc is
    port (
        clk           : in  std_logic;                      
        rst           : in  std_logic;                      
    -- ir e pc
        opcode_in     : in  unsigned(3 downto 0);          -- opcode [16:13] 
        pc_atual_in   : in  unsigned(16 downto 0);          -- pc
        const_5bit_in : in  unsigned(4 downto 0);          -- constante [4:0] 
        const_13bit_in: in  unsigned(12 downto 0);         -- endereço [12:0] pro jump 
--saidas
        pc_wr_en_out  : out std_logic;                      -- escrita no PC
        ir_wr_en_out  : out std_logic;                      -- escrita no IR
        reg_wr_en_out : out std_logic;                      -- escrita no banco
        ula_chave_out : out std_logic_vector(1 downto 0);   -- operação da ula
        sel_mux_ula_b_out : out std_logic;                  -- entrada B da ula
        sel_mux_reg_wr_out: out std_logic;                 -- dado a escrever no banco, 0 ula 1 banco
        pc_in_out     : out unsigned(16 downto 0)           -- próximo pc
    );
end entity uc;

architecture a_uc of uc is

  component maq_estados is
    port ( 
        clk,rst: in std_logic;
        estado: out unsigned(1 downto 0)
    );
  end component;

  signal s_estado_atual: unsigned(1 downto 0);

begin

state_instance: maq_estados
  port map (
          clk => clk,
          rst => rst,
          estado => s_estado_atual
    );

  ir_wr_en_out <= '1' when s_estado_atual = "00" else '0'; --fetch

  pc_wr_en_out <= '1' when s_estado_atual = "01" else '0'; --decode

  pc_in_out <= ("0000" & const_13bit_in) when (s_estado_atual = "01" and opcode_in = "1111") else --jump
               (pc_atual_in + 1) when (s_estado_atual = "01") else --pc + 1
               pc_atual_in; --mantem

  --controle do banco
  reg_wr_en_out <= '1' when (s_estado_atual = "10") and
                   (opcode_in = "0001" or --add 
                    opcode_in = "0010" or --sub 
                    opcode_in = "1000" or --addi
                    opcode_in = "1001") --subi
                  else '0';
    
    --controele da ull 
    ula_chave_out <= "00" when (s_estado_atual = "10") and (opcode_in = "0001" or opcode_in = "1000") else --add e addi 
                     "01" when (s_estado_atual = "10") and (opcode_in = "0010" or opcode_in = "1001") else --sub e subi
                     "00"; -- nop, jump etc 
                   
    --mux da ula
    sel_mux_ula_b_out <= '1' when (s_estado_atual = "10") and 
                         (opcode_in = "1000" or -- addi
                         opcode_in = "1001") -- subi
                       else '0'; --por padrao pega do registrador

    --mux do banco 
      sel_mux_reg_wr_out <= '1' when (s_estado_atual = "10") and
                            (opcode_in = "1000") --addi
                          else '0'; --saida da ula

end architecture a_uc;
