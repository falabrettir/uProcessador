library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(16 downto 0)
   );
end entity;

architecture a_rom of rom is

   type mem is array (0 to 127) of unsigned(16 downto 0);
   constant conteudo_rom : mem := (
      
-- ===============================================================
      -- 1. INICIALIZAÇÃO (R1=79, R4=33, R7=0)
      -- ===============================================================
      0  => "00100001000100010", -- CLR R1
      1  => "10000001000101111", -- ADDI R1, 15
      2  => "10000001000101111", -- ADDI R1, 15
      3  => "10000001000101111", -- ADDI R1, 15
      4  => "10000001000101111", -- ADDI R1, 15
      5  => "10000001000101111", -- ADDI R1, 15
      6  => "10000001000100100", -- ADDI R1, 4 (R1=79)

      7  => "00100010001000100", -- CLR R2
      8  => "10000010001001111", -- ADDI R2, 15
      9  => "10000010001001111", -- ADDI R2, 15
      10 => "10000010001000011", -- ADDI R2, 3
      11 => "11100100001000000", -- MOV R4, R2 (R4=33)

      12 => "00100111011101110", -- CLR R7 (Zero)

      -- ===============================================================
      -- 2. PREENCHIMENTO RAM (0..32)
      -- ===============================================================
      13 => "00100010001000100", -- CLR R2 (i=0)

      -- LOOP FILL (End 14)
      14 => "11100011000100000", -- MOV R3, R1 (Base)
      15 => "00010011001000000", -- ADD R3, R2 (Base + i)
      
      -- SW CORRIGIDO: Dado R2(12-9), Addr R3(8-5)
      -- Bin: 1011 0010 0011 00000
      16 => "10110010001100000", -- SW R2, (R3)
      
      17 => "10000010001000001", -- ADDI R2, 1
      18 => "00110010010000000", -- CMPR R2, R4
      19 => "11011111111111010", -- BLO -6

      -- 2B. LIMPEZA DO 0 e 1 (End 79 e 80)
      -- SW R7(Zero), (R1=79) -> Dado R7(12-9), Addr R1(8-5)
      20 => "10110111000100000", 
      
      21 => "11100011000100000", -- MOV R3, R1
      22 => "10000011001100001", -- ADDI R3, 1 (80)
      -- SW R7, (R3) -> Dado R7, Addr R3
      23 => "10110111001100000", 

      -- ===============================================================
      -- 3. CRIVO DO 2
      -- ===============================================================
      24 => "00100101010100101", -- CLR R5
      25 => "10000101010100010", -- ADDI R5, 2
      26 => "11100110010100000", -- MOV R6, R5

      -- LOOP 2 (End 27)
      27 => "00010110010100000", -- ADD R6, R5
      28 => "00110110010000000", -- CMPR R6, R4
      29 => "11010000000000001", -- BLO +1
      30 => "11110000000100101", -- JMP 37 (Sai)

      -- WRITE (End 31)
      31 => "11100011000100000", -- MOV R3, R1
      32 => "00010011011000000", -- ADD R3, R6
      -- SW R7, (R3) -> Dado R7(12-9), Addr R3(8-5)
      33 => "10110111001100000", 
      34 => "11110000000011011", -- JMP 27

      -- ===============================================================
      -- 4. CRIVO DO 3
      -- ===============================================================
      35 => "00000000000000000", -- Padding
      36 => "00000000000000000",

      37 => "00100101010100101", -- CLR R5
      38 => "10000101010100011", -- ADDI R5, 3
      39 => "11100110010100000", -- MOV R6, R5

      -- LOOP 3 (End 40)
      40 => "00010110010100000", 
      41 => "00110110010000000",
      42 => "11010000000000001",
      43 => "11110000000110010", -- JMP 50

      44 => "11100011000100000",
      45 => "00010011011000000",
      -- SW R7, (R3)
      46 => "10110111001100000",
      47 => "11110000000101000", -- JMP 40

      -- ===============================================================
      -- 5. CRIVO DO 5
      -- ===============================================================
      48 => "00000000000000000",
      49 => "00000000000000000",

      50 => "00100101010100101", -- CLR R5
      51 => "10000101010100101", -- ADDI R5, 5
      52 => "11100110010100000", -- MOV R6, R5

      -- LOOP 5 (End 53)
      53 => "00010110010100000",
      54 => "00110110010000000",
      55 => "11010000000000001",
      56 => "11110000000111101", -- JMP 61

      57 => "11100011000100000",
      58 => "00010011011000000",
      -- SW R7, (R3)
      59 => "10110111001100000",
      60 => "11110000000110101", -- JMP 53

      -- ===============================================================
      -- 6. LEITURA FINAL
      -- ===============================================================
      61 => "00100101010100000", -- CLR R5 (Comparador de inteiros)
      62 => "00101000100000000", -- CLR R8 (Pino de saída) 
      
      63 => "00100010001000000", -- CLR R2

      -- READ LOOP (End 64)
      64 => "10000010001000001", -- ADDI R2, 1 
      
      65 => "11100011000100000", -- MOV R3, R1
      66 => "00010011001000000", -- ADD R3, R2
      
      -- LW R7, (R3) -> Dest R7(12-9), Addr R3(8-5)
      -- Hardware LW lê bits 8-5 para endereço.
      67 => "01110111001100000", 
            
      68 => "00100101010100000", -- CLR R5 (Zera R5 antes de acumular)
      69 => "01000101011100000", --OR R5, R7 (Acumula em R5)
      
      70 => "00110000010100000", --CMPR R0, R5 (FLAGS: R0-R5)

      71 => "11010000000000100", --BLO +4 (SE R5 > 0, manda pra saida (PC=75))
        
      72 => "00110010010000000", -- CMPR R2, R4 (FLAGS: R2-R4)

      73 => "11010000000000001", -- BLO +1 (se R2 < R4, continua leitura)
      
      74 => "11110000001001010", -- HALT (CABOU.)

      75 => "11011111111110100", -- BLO -12 (loop de leitura em PC=64)

      76 => "11101000011100000", --MOV R8, R7 (Saída)
      77 => "11110000001000000", --JMP 64 (volta para o loop de leitura)

      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture a_rom;
