library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(16 downto 0)
   );
end entity;

architecture a_rom of rom is

   type mem is array (0 to 127) of unsigned(16 downto 0);
   constant conteudo_rom : mem := (
      
      0  => "00100001000100010", -- CLR R1
      1  => "10000001000101111", -- ADDI R1, 15
      2  => "10000001000101111", -- ADDI R1, 15
      3  => "10000001000101111", -- ADDI R1, 15
      4  => "10000001000101111", -- ADDI R1, 15
      5  => "10000001000101111", -- ADDI R1, 15
      6  => "10000001000100100", -- ADDI R1, 4 (R1=79)

      7  => "00100010001000100", -- CLR R2
      8  => "10000010001001111", -- ADDI R2, 15
      9  => "10000010001001111", -- ADDI R2, 15
      10 => "10000010001000011", -- ADDI R2, 3
      11 => "11100100001000000", -- MOV R4, R2 (R4=33)
      
      12 => "00100111011101110", -- CLR R7 (Zero)

      -- 2. PREENCHIMENTO RAM (0..32)
      13 => "00100010001000100", -- CLR R2 (i=0)

      -- LOOP FILL (End 14)
      14 => "11100011000100000", -- MOV R3, R1 (Base)
      15 => "00010011001000000", -- ADD R3, R2 (Base + i)
      
      -- Bin: 1011 0010 0011 00000
      16 => "10110010001100000", -- SW R2, (R3)
      
      17 => "10000010001000001", -- ADDI R2, 1
      18 => "00110010010000000", -- CMPR R2, R4
      19 => "11011111111111010", -- BLO -6

      -- 2B. LIMPEZA DO 0 e 1 (End 79 e 80)
      -- SW R7(Zero), (R1=79) -> Dado R7(12-9), Addr R1(8-5)
      20 => "10110111000100000", 
      
      21 => "11100011000100000", -- MOV R3, R1
      22 => "10000011001100001", -- ADDI R3, 1 (80)
      -- SW R7, (R3) -> Dado R7, Addr R3
      23 => "10110111001100000", 

      24 => "00100010001000100", -- CLR R2
      25 => "10000010001001111", -- ADDI R2, 15
      26 => "10000010001001111", -- ADDI R2, 15
      27 => "10000010001000001", -- ADDI R2, 1
      -- máscara de bits
      -- 3. CRIVO DO 2
      28 => "00100101010100101", -- CLR R5
      29 => "10000101010100010", -- ADDI R5, 2
      30 => "11100110010100000", -- MOV R6, R5
                                 -- LOOP 2 START
      -- 1. Incrementa
      31 => "00010110010100000", -- ADD R6, R5
      
      -- Grava Zero na posição RAM[79 + R6]
      32 => "11100011000100000", -- MOV R3, R1 (Base 79)
      33 => "00010011011000000", -- ADD R3, R6 (Endereço Absoluto)
      34 => "10110111001100000", -- SW R7, (R3) (Escreve 0)
      
      35 => "11101000011000000", -- MOV R8, R6
      36 => "01001000001000000", -- OR  R8, R2 
      37 => "00111000001000000", -- CMPR R8, R2
      
      -- 4. Decisão
      -- Se Z=0 (Deu 63), sai. 
      -- BNE +1 
      38 => "11000000000000001", -- BNE +1 (Vai para 40)

      -- 5. Volta
      -- JMP para 31 (ADD R6, R5)
      39 => "11110000000011111", -- JMP 31

      -- 4. CRIVO DO 3
      -- Inicialização (R5=3, R6=3)
      40 => "00100101010100101", -- CLR R5
      41 => "10000101010100011", -- ADDI R5, 3
      42 => "11100110010100000", -- MOV R6, R5

      -- LOOP 3 START (Endereço 43)
      -- 1. Incrementa (R6 = 6, 9, 12...)
      43 => "00010110010100000", -- ADD R6, R5
      
      -- 2. Escrita na Memória
      44 => "11100011000100000", -- MOV R3, R1 (Base 79)
      45 => "00010011011000000", -- ADD R3, R6 (Endereço = 79 + R6)
      46 => "10110111001100000", -- SW R7, (R3) (Escreve 0)

      -- 3. Verificação com Máscara OR (R2 ainda tem 31)
      47 => "11101000011000000", -- MOV R8, R6
      48 => "01001000001000000", -- OR  R8, R2 (R8 = R6 OR 31)
      49 => "00111000001000000", -- CMPR R8, R2 (Deu 31?)
      
      -- Pula para linha 52
      50 => "11000000000000001", -- BNE +1 

      -- JMP para 43 (ADD R6, R5)
      51 => "11110000000101011", -- JMP 43
      
      52 => "00000000000000000", -- NOP 


      -- 5. CRIVO DO 5
      -- Inicialização (R5=5, R6=5)
      53 => "00100101010100101", -- CLR R5
      54 => "10000101010100101", -- ADDI R5, 5
      55 => "11100110010100000", -- MOV R6, R5

      -- LOOP 5 START (Endereço 56)
      -- 1. Incrementa (R6 = 10, 15, 20...)
      56 => "00010110010100000", -- ADD R6, R5

      -- 2. Escrita na Memória
      57 => "11100011000100000", -- MOV R3, R1 (Base 79)
      58 => "00010011011000000", -- ADD R3, R6 (Endereço = 79 + R6)
      59 => "10110111001100000", -- SW R7, (R3)

      -- 3. Verificação com Máscara OR
      60 => "11101000011000000", -- MOV R8, R6
      61 => "01001000001000000", -- OR  R8, R2
      62 => "00111000001000000", -- CMPR R8, R2
      
      -- 4. Decisão
      -- Se Z=0, sai. BNE +1 (Pula o JMP). Vai para 65.
      63 => "11000000000000001", -- BNE +1

      -- 5. Volta
      -- JMP para 56 (ADD R6, R5)
      64 => "11110000000111000", -- JMP 56 

      65 => "00000000000000000", -- NOP / Padding
      -- leitura
      66 => "00100101010100000", -- CLR R5 (Comparador de inteiros)
      67 => "00101000100000000", -- CLR R8 (Pino de saída) 
      
      68 => "00100010001000000", -- CLR R2

      -- READ LOOP (End 64)
      69 => "10000010001000001", -- ADDI R2, 1 
      
      70 => "11100011000100000", -- MOV R3, R1
      71 => "00010011001000000", -- ADD R3, R2
      
      -- LW R7, (R3) -> Dest R7(12-9), Addr R3(8-5)
      -- Hardware LW lê bits 8-5 para endereço.
      72 => "01110111001100000", 
            
      73 => "00100101010100000", -- CLR R5 (Zera R5 antes de acumular)
      74 => "01000101011100000", --OR R5, R7 (Acumula em R5)
      
      75 => "00110000010100000", --CMPR R0, R5 (FLAGS: R0-R5)

      76 => "11010000000000100", --BLO +4 (SE R5 > 0, manda pra saida (PC=75))
        
      77 => "00110010010000000", -- CMPR R2, R4 (FLAGS: R2-R4)

      78 => "11010000000000001", -- BLO +1 (se R2 < R4, continua leitura)
      
      79 => "11110000001001010", -- HALT (CABOU.)

      80 => "11011111111110100", -- BLO -12 (loop de leitura em PC=64)

      81 => "11101000011100000", --MOV R8, R7 (Saída)
      82 => "11110000001000000", --JMP 64 (volta para o loop de leitura)

      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture a_rom;
